* exp3.cir
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=55                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     Vdd     0       2.5
***********************************************************************
* Define Subcircuits
***********************************************************************
.subckt front_inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=32u
m2      Out In Vdd Vdd  cmosp l=0.25u w=64u
.ends

.subckt end_inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=2u
m2      Out In Vdd Vdd  cmosp l=0.25u w=4u
.ends
***********************************************************************
* Stimulus
***********************************************************************
* Format of pulse input:
*Vin     In      0       PULSE(0 2.5 1n 0.1n 0.1n 4n 10n)
*V1       In      0       PWL(0n 0 0.1n 1)
V1       In      0       PWL(0n 0 1n 0 2n 2.5)
***********************************************************************

* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here
**1-1段**
*R1 In a 100
*C1  a 0 100p

**1-2段**
*R1 In a 100
*R2  a b 100
*C1  a 0 100p
*C2  b 0 100p

*1-3段*
*R1 In a 100
*R2  a b 100
*R3  b c 100
*C1  a 0 100p
*C2  b 0 100p
*C3  c 0 100p

*2*
*R=0.08/□, C=0.32fF/um, 2mm 0.5um
*0.08 * 2 / 0.5 => 0.32 で考える
*コンデンサについては 0.32 * 2000 = 640fFを分割

x0 In a Vdd front_inv
**pi 1**
*C1 a 0 320f
*R1 a b 0.32
*C2 b 0 320f

**T 1 **
R1 a b 0.16
C1 b 0 640f
R2 b c 0.16

x1 c Out Vdd end_inv
Ce Out 0 12f
*******************************************


.tran 0.001ns 12ns
.plot TRAN V(In) V(a) V(b) V(c) V(Out) V(d) V(e)
***********************************************************************
* End of Deck
***********************************************************************
.end
