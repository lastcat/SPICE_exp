* sample.cir
* ゲートテスト用の回路
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=55                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     Vdd     0       2.5
***********************************************************************
* Define Subcircuits
***********************************************************************
.subckt inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=2u
m2      Out In Vdd Vdd  cmosp l=0.25u w=4u
.ends
.subckt inva In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=4u
m2      Out In Vdd Vdd  cmosp l=0.25u w=8u
.ends
.subckt invb In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=16u
m2      Out In Vdd Vdd  cmosp l=0.25u w=32u
.ends
.subckt invc In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=64u
m2      Out In Vdd Vdd  cmosp l=0.25u w=128u
.ends

*2入力NAND
.subckt t_nand in_a in_b Out Vdd
*m1   　　Drain Gate Source 基盤? cmons(n/p) l=0.25u w=3u
m1        Vdd in_a Out Vdd cmosp l=0.25u w=6u
m2        Out   in_a b 0   cmosn l=0.25u w=6u
m3        b   in_b 0 0   cmosn l=0.25u w=6u
m4        Vdd in_b Out Vdd cmosp l=0.25u w=6u
.ends

*2入力NOR
.subckt t_nor in_a in_b Out Vdd
m1    Vdd in_a a Vdd cmosp l=0.25u w=6u
m2    a   in_b Out Vdd cmosp l=0.25u w=6u
m3    Out   in_b 0 0   cmosn l=0.25u w=6u
m4    Out   in_a 0 0   cmosn l=0.25u w=6u
.ends

*4入力NAND
.subckt f_nand in_a in_b in_c in_d Out Vdd
m1    Vdd in_a Out Vdd cmosp l=0.25u w=6u
m2    Out in_a a   0   cmosn l=0.25u w=6u
m3    a   in_b b   0   cmosn l=0.25u w=6u
m4    b   in_c c   0   cmosn l=0.25u w=6u
m5    c   in_d 0   0   cmosn l=0.25u w=6u
m6    Vdd in_b Out Vdd cmosp l=0.25u w=6u
m7    vdd in_c Out Vdd cmosp l=0.25u w=6u
m8    Vdd in_d Out Vdd cmosp l=0.25u w=6u
.ends

*4入力NOR
.subckt f_nand in_a in_b in_c in_d Out Vdd
m1    0 in_a Out 0 cmosn l=0.25u w=6u
m2    Out in_a a   Vdd   cmosp l=0.25u w=6u
m3    a   in_b b   Vdd   cmosp l=0.25u w=6u
m4    b   in_c c   Vdd   cmosp l=0.25u w=6u
m5    c   in_d Vdd   Vdd   cmosp l=0.25u w=6u
m6    0 in_b Out 0 cmosn l=0.25u w=6u
m7    0 in_c Out 0 cmosn l=0.25u w=6u
m8    0 in_d Out 0 cmosn l=0.25u w=6u
.ends

*これで試して今日のこれは終わり まあ少しずつ勉強していってもいいかな
***********************************************************************
* Stimulus
***********************************************************************
* Format of pulse input:
* pulse v_initial v_final t_delay t_rise t_fall t_pulsewidth t_period
Vin     in_one      0       PULSE(0 2.5 1ns 0.1ns 0.1ns 4ns 10ns)
*Vin     in_one      0       1
V1      in_two      0       0
***********************************************************************
* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here

x1      in_one    in_two    Out     Vdd t_nor
*x2      a       b       Vdd     inva
*r1      b       c       1k
*c1      c       0       100f
*r2      c       Out     1k
*x4      Out     d       Vdd     invb
*x5      d       e       Vdd     invc
.tran .001ns 12ns
.plot TRAN V(In) V(a) V(b) V(c) V(Out) V(d) V(e)
***********************************************************************
* End of Deck
***********************************************************************
.end
