* exp4_1.cir
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=27                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     Vdd     0       2.5
***********************************************************************
* Define Subcircuits
***********************************************************************
.subckt inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=2u
m2      Out In Vdd Vdd  cmosp l=0.25u w=4u
.ends

***********************************************************************
* Stimulus
***********************************************************************
* Format of pulse input:
* pulse v_initial v_final t_delay t_rise t_fall t_pulsewidth t_period
Vin     In      0       PWL(0n 2.5 1.0n 2.5 3n 0 6.0n 0 8n 2.5 10.0n 2.5)
***********************************************************************
* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here

x1 in Out Vdd inv
c1 Out 0 64f
*0.1n =>  1.532285e-05
*1n => 2.393863e-05
*2n => 3.615765e-0
*あとは計算*

.tran .001ns 12ns
.plot TRAN V(In) V(a) V(b) V(c) V(Out) V(d) V(e)
***********************************************************************
* End of Deck
***********************************************************************
.end
