* exp3.cir
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=55                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     Vdd     0       2.5
***********************************************************************
* Define Subcircuits
***********************************************************************
.subckt front_inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=32u
m2      Out In Vdd Vdd  cmosp l=0.25u w=64u
.ends

.subckt end_inv In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=2u
m2      Out In Vdd Vdd  cmosp l=0.25u w=4u
.ends

***********************************************************************
* Stimulus
***********************************************************************
* Format of pulse input:
*3-1用電流*
*V1       In      0       PWL(0n 0 0.1n 1)
*3-2用電流*
Vin     In      0       PULSE(0 2.5 1n 0.1n 0.1n 1n 3n)

*V1       In      0       PWL(0n 0 1n 0 2n 2.5 3n 2.5 4n 0)
***********************************************************************

* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here
**3-1**
**1-1段**
*比較用の一段回路　Rの値は適宜修正
*R1 In a 600
*C1  a 0 100p

**1-2段**
*R1 In a 100
*R2  a b 100
*C1  a 0 100p
*C2  b 0 100p

*1-3段*
*R1 In a 100
*R2  a b 100
*R3  b c 100
*C1  a 0 100p
*C2  b 0 100p
*C3  c 0 100p

*3-2*
*R=0.08/□, C=0.32fF/um, 2mm 0.5um
*0.08 * 2 / 0.5 * 1000 => 320
*コンデンサについては 0.32 * 2000 = 640fFを分割
*PULSEの上り(1.25v)　1.05e-09 下り(1.25v) 2.15e-09

**手前のインバーター**
x0 In a Vdd front_inv

**pi_1** 
*C1 a 0 320f
*R1 a b 320
*C2 b 0 320f

**pi_2** 
*C1 a 0 160f
*R1 a b 160
*C2 b 0 320f
*R2 b c 160
*C3 c 0 160f

**l_1**
*R1 a b 320
*C1 b 0 640f 

**l_4**
R1 a b 80
C1 b 0 160f
R2 b c 80
C2 c 0 160f
R3 c d 80
C3 d 0 160f
R4 d e 80
C4 e 0 160f

**t_1 **
*R1 a b 160
*C1 b 0 640f
*R2 b c 160

**t_2 **
*R1 a b 80
*C1 b 0 320f
*R2 b c 160
*C2 c 0 320f
*R3 c d 80


x1 e Out Vdd end_inv
C100 Out 0 12f
*******************************************


.tran 0.001ns 10ns
.plot TRAN V(In) V(a) V(b) V(c) V(Out) V(d) V(e)
***********************************************************************
* End of Deck
***********************************************************************
.end
